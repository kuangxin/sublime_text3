module test (
    input  logic                    i_en            ,
    output logic [pq_symbols*4-1:0] o_all_symbols_4b,
    input  logic                    i_en2
);
endmodule