module t #(
    aa = 1,

    bb = 2
) (
    input  logic a,

    output logic b,

    output logic c
);
endmodule